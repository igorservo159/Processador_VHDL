library ieee;
use ieee.std_logic_1164.all;

entity processor is
	Port(
		clk_pro: in std_logic;
	);
end processor;

architecture behav of processor is
	component datapath is
		Port(
			clk_dp: in std_logic;
	
			D_addr: in std_logic_vector(7 downto 0);
			D_rd, D_wr: in std_logic;
	
			RF_W_data: in std_logic_vector(15 downto 0);
			RF_s1, RF_s0: in std_logic;
			
			RF_W_addr: in std_logic_vector(3 downto 0);
			RF_W_wr: in std_logic;
			
			RF_Rp_addr: in std_logic_vector(3 downto 0);
			RF_Rp_rd: in std_logic;
	
			RF_Rq_addr: in std_logic_vector(3 downto 0);
			RF_Rq_rd: in std_logic;
	
			RF_Rp_zero: out std_logic;
			
			ALU_s1, ALU_s0: in std_logic);
	end component;
	
	component control_unit is
		Port(
			clk_ctl_un, RP_zero_ctl_un: in std_logic;
			
			alu_s0_ctl_un, alu_s1_ctl_un: out std_logic;
			
			D_wr_ctl_un, D_rd_ctl_un: out std_logic;
			D_addr_ctl_un: out std_logic_vector(8 downto 0);
			
			W_addr_ctl_un, Rp_addr_ctl_un, Rq_addr_ctl_un: out std_logic_vector(4 downto 0);
			Rp_rd_ctl_un, Rq_rd_ctl_un, W_wr_ctl_un, RF_s0_ctl_un, RF_s1_ctl_un: out std_logic;
			W_data_ctl_un: out std_logic_vector(15 downto 0));
	end component;
	
	signal RP_zero_pro: std_logic;
	signal alu_s0_pro, alu_s1_pro:std_logic;
	signal D_wr_pro, D_rd_pro:std_logic;
	signal D_addr_pro:std_logic_vector(8 downto 0);
	signal W_addr_pro, Rp_addr_pro, Rq_addr_pro: std_logic_vector(4 downto 0);
	signal Rp_rd_pro, Rq_rd_pro, W_wr_pro, RF_s0_pro, RF_s1_pro: std_logic;
	signal W_data_pro: std_logic_vector(15 downto 0);

	begin
		u1: datapath port map(clk_dp=>clk_pro, D_addr=>D_addr_pro, D_rd=>D_rd_pro, D_wr=>D_wr_pro,
							  RF_W_data=>W_data_pro, RF_W_addr,
							  RF_W_wr, RF_s1=>RF_s0_pro, RF_s0=> RF_s1_pro,
							  RF_Rp_addr=>Rp_addr_pro, RF_Rp_rd=>Rp_rd_pro, RF_Rp_zero=>RP_zero_pro,
							  ALU_s1=>alu_s1_pro, ALU_s0=>alu_s0_pro);

		u2: control_unit port map(clk_ctl_un=>clk_pro, RP_zero_ctl_un=>RP_zero_pro,
								  alu_s0_ctl_un=>alu_s0_pro, alu_s1_ctl_un=>alu_s1_pro,
								  D_wr_ctl_un=>D_wr_pro, D_rd_ctl_un=>D_rd_pro, D_addr_ctl_un=>D_addr_pro,
								  W_addr_ctl_un=>W_addr_pro, Rp_addr_ctl_un=>Rp_addr_pro,
								  Rq_addr_ctl_un=>Rq_addr_pro, Rp_rd_ctl_un=>Rp_rd_pro,
								  Rq_rd_ctl_un=>Rq_rd_pro, W_wr_ctl_un=>W_wr_pro,
								  RF_s0_ctl_un=>RF_s0_pro, RF_s1_ctl_un=>RF_s1_pro, W_data_ctl_un=>W_data_pro);
end behav;